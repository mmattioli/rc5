--
-- Written by Michael Mattioli
--
--
-- Description: Key expansion module.
--
