--
-- Written by Michael Mattioli
--
--
-- Description: RC5 decryption module.
--
