--
-- Written by Michael Mattioli
--
--
-- Description: RC5 encryption module.
--
